grammar silver:driver;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Driver\nmenu_title: Driver\nmenu_weight: 100\n---"
@}

