grammar edu:umn:cs:melt:tutorial:expr:host_op_overloading ;

-- This file defines the new addition operator that 
-- supports operator overloading.

import edu:umn:cs:melt:tutorial:expr:terminals ;
import edu:umn:cs:melt:tutorial:expr:abstractsyntax ;
import edu:umn:cs:melt:tutorial:expr:concretesyntax ;



-- Concrete Syntax --
---------------------

-- This is the new concrete syntax for addition and it replaces
-- 'add' in expr:concretesyntax.  This new production creates 
-- an AST using the new add_overload production.  

concrete production add_overload_c
sum::Expr_c ::= e::Expr_c  op::Plus_t  t::Expr_c
{
 sum.pp = e.pp ++ " " ++ op.lexeme ++ " " ++ t.pp ;
 sum.ast_Expr = add_overload(e.ast_Expr, op, t.ast_Expr );
}


-- Abstract Syntax --
---------------------

-- This production provides the "extension point" or "hook" that
-- language extensions can use to overload the addition operator.

-- This is done by using a production attriubte 'overloads' that is
-- populated by language extensions (and the aspect production furter
-- below).   Aspect productions on add_overload will typically examine
-- the types (typerep attributes) on the two children to see if they
-- are the types of interest, and if so, the aspect production wil create
-- a new AST that the add_overload production should forward to.

-- If the number of trees in 'overloads' is not 1, an error message is
-- generated by forwarding to the error_Expr production.

abstract production add_overload
sum::Expr ::= l::Expr  op::Plus_t  r::Expr
{
 sum.pp = "(" ++ l.pp ++ " " ++ op.lexeme ++ " " ++ r.pp ++ ")";

 production attribute overloads :: [ Expr ] with ++ ;
 overloads := [ ] ;

 forwards to
   if   length(overloads) == 1
   then head(overloads)
   else
   if   length(overloads) == 0
   then error_Expr (
          op.line, op.column,
          "Addition not supported on types " ++
          l.typerep.pp ++ " and " ++ r.typerep.pp ) 
   else error_Expr (
          op.line, op.column,
          "Addition implemented in multiple ways on types " ++
          l.typerep.pp ++ " and " ++ r.typerep.pp ) ;
}



-- Overload + for integer addition.  Thus, integer expressions
-- that were valid in the orignial (expr:host) language are also
-- valid in this language that supports overloading.

aspect production add_overload
sum::Expr ::= l::Expr op::Plus_t  r::Expr
{
 overloads <- if   equal_types(l.typerep, intType()) &&
                   equal_types(r.typerep, intType())
              then [ add(l,op,r) ] 
              else [ ] ;
}



