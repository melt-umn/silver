grammar silver:compiler:extension:abella_compilation;

imports silver:compiler:definition:core;
imports silver:compiler:definition:env;

imports silver:compiler:driver:util;

imports silver:compiler:extension:abella_compilation:encoding;
imports silver:compiler:extension:abella_compilation:abella;
imports silver:compiler:extension:abella_compilation:parsing_thms;

