grammar copper_features;

imports silver:testing ;
imports lib:extcore ;

import copper_features:test_layout;

mainTestSuite copper_tests ;

{- Needed: 
layout tests
precedence / associativity tests
lexer classes & dominates submits tests
production precedence / operator tests
-}
