grammar edu:umn:cs:melt:tutorial:expr:abstractsyntax ;

-- Operator overloading is not supported in the original
-- version of the tutorial:expr language. 

-- It is added in the grammars
--  expr:host:op_overloading
--  expr:exts:float
--  expr:composed:expr_float

-- These are provided to illustrate how operator overloading works in
-- the extensible Java specifications in ableJ and in other language
-- specifications.

-- Since this expression grammar is used for tutorials, we decided to
-- keep the host language as simple as possible and that led us to
-- leave operator overloading out of the host language.
