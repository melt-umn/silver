

import silver_features:defs:subdefs as c;


synthesized attribute newattr :: c:Bar;

