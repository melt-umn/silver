grammar silver:langutil;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Language Utilities\nmenu_title: Lang Util\nmenu_weight: 100\n---"
@}

