grammar silver_features:cond:d;

exports silver_features:cond:e with silver_features:cond:d;

global bVal :: Integer = 5;
