grammar silver:definition:concrete_syntax;

imports silver:definition:core;
imports silver:definition:type:syntax;

imports silver:definition:env;
imports silver:definition:type;

imports silver:definition:concrete_syntax:ast;

option silver:modification:copper;

exports silver:definition:concrete_syntax:ast:env_parser with silver:definition:env:env_parser;
