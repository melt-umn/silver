grammar lib:lsp:document;

imports lib:lsp:json;
imports lib:lsp;
