grammar silver:core;

data Unit = unit;
derive Eq, Ord on Unit;
