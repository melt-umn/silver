grammar silver;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Silver\nmenu_title: Silver\nmenu_weight: 100\n---"
@}

