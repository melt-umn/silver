grammar silver:modification:propagatedattribs;

imports silver:definition:core;
imports silver:definition:type:syntax;

imports silver:definition:env;
imports silver:definition:type;

import silver:util;