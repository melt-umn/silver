
monoid attribute defs::[String] with [], ++;
monoid attribute freeVars::[String] with [], ++;

propagate defs on MStmt;
propagate freeVars on MExpr;

nonterminal MStmt with defs, freeVars;
nonterminal MExpr with freeVars;

abstract production seqMStmt
top::MStmt ::= s1::MStmt s2::MStmt
{
  top.freeVars := s1.freeVars ++ removeAllBy(stringEq, s1.defs, s2.freeVars);
}

abstract production assignMStmt
top::MStmt ::= a::String e::MExpr
{
  propagate freeVars;
  top.defs <- [a];
}

abstract production addMExpr
top::MExpr ::= e1::MExpr e2::MExpr
{}

abstract production varMExpr
top::MExpr ::= a::String
{
  top.freeVars <- [a];
}

global testMStmt::MStmt =
  seqMStmt(
    assignMStmt("a", addMExpr(varMExpr("b"), varMExpr("c"))),
    assignMStmt("d", varMExpr("a")));

equalityTest(testMStmt.defs, ["a", "d"], [String], silver_tests);
equalityTest(testMStmt.freeVars, ["b", "c"], [String], silver_tests);
