grammar silver:extension:bidirtransform;
