grammar silver:core;

nonterminal IOMonad<a> with stateIn<IO>, stateOut<IO>, stateVal<a>;

abstract production bindIO
top::IOMonad<b> ::= st::IOMonad<a> fn::(IOMonad<b> ::= a)
{
  st.stateIn = top.stateIn;
  local newState::IOMonad<b> = fn(st.stateVal);
  newState.stateIn = st.stateOut;
  local stateOut::IO = newState.stateOut;
  local stateVal::b = newState.stateVal;
  
  -- Using unsafeTrace here to demand st is evaluated before evaluating fn
  top.stateOut = unsafeTrace(stateOut, st.stateOut);
  top.stateVal = unsafeTrace(stateVal, st.stateOut);
}

abstract production returnIO
top::IOMonad<a> ::= x::a
{
  top.stateOut = top.stateIn;
  top.stateVal = x;
}

instance Functor IOMonad {
  map = liftM1;
}

instance Apply IOMonad {
  ap = apM;
}

instance Applicative IOMonad {
  pure = returnIO;
}

instance Bind IOMonad {
  bind = bindIO;
}

instance Monad IOMonad {}

function runIO
IO ::= st::IOMonad<a> ioIn::IO
{
  return evalIO(st, ioIn).io;
}

function evalIO
IOVal<a> ::= st::IOMonad<a> ioIn::IO
{
  st.stateIn = ioIn;
  return ioval(st.stateOut, st.stateVal);
}

function unsafeEvalIO
a ::= st::IOMonad<a>
{
  return evalIO(st, unsafeIO()).iovalue;
}

-- Monadic IO wrappers
abstract production wrapIOToken
top::IOMonad<Unit> ::= f::(IO ::= IO)
{
  top.stateOut = f(top.stateIn);
  top.stateVal = unit();
}

abstract production wrapIOVal
top::IOMonad<a> ::= f::(IOVal<a> ::= IO)
{
  local res::IOVal<a> = f(top.stateIn);
  top.stateOut = res.io;
  top.stateVal = res.iovalue;
}

abstract production printM
top::IOMonad<Unit> ::= s::String
{ forwards to wrapIOToken(print(s, _)); }

abstract production readLineStdinM
top::IOMonad<String> ::=
{ forwards to wrapIOVal(readLineStdin); }

-- Having a polymorphic return type lets us write code like:
--
--   if !null(errs) {
--     printM(showErrs(errs));
--     exitM(1);
--   } else {
--     return value;
--   }
abstract production exitM
top::IOMonad<a> ::= val::Integer
{
  top.stateOut = exit(val, top.stateIn);
  top.stateVal = error("stateOut should've been evaluated first?");
}

abstract production mkdirM
top::IOMonad<Boolean> ::= s::String
{ forwards to wrapIOVal(mkdir(s, _)); }

abstract production systemM
top::IOMonad<Integer> ::= s::String
{ forwards to wrapIOVal(system(s, _)); }

abstract production writeFileM
top::IOMonad<Unit> ::= file::String contents::String
{ forwards to wrapIOToken(writeFile(file, contents, _)); }

abstract production appendFileM
top::IOMonad<Unit> ::= file::String contents::String
{ forwards to wrapIOToken(appendFile(file, contents, _)); }

abstract production fileTimeM
top::IOMonad<Integer> ::= s::String
{ forwards to wrapIOVal(fileTime(s, _)); }

abstract production isFileM
top::IOMonad<Boolean> ::= s::String
{ forwards to wrapIOVal(isFile(s, _)); }

abstract production isDirectoryM
top::IOMonad<Boolean> ::= s::String
{ forwards to wrapIOVal(isDirectory(s, _)); }

abstract production readFileM
top::IOMonad<String> ::= s::String
{ forwards to wrapIOVal(readFile(s, _)); }

abstract production cwdM
top::IOMonad<String> ::= 
{ forwards to wrapIOVal(cwd); }

abstract production envVarM
top::IOMonad<String> ::= s::String
{ forwards to wrapIOVal(envVar(s, _)); }

abstract production listContentsM
top::IOMonad<[String]> ::= s::String
{ forwards to wrapIOVal(listContents(s, _)); }

abstract production deleteFileM
top::IOMonad<Boolean> ::= s::String
{ forwards to wrapIOVal(deleteFile(s, _)); }

abstract production deleteTreeM
top::IOMonad<Unit> ::= s::String
{ forwards to wrapIOToken(deleteTree(s, _)); }

abstract production copyFileM
top::IOMonad<Unit> ::= src::String dst::String
{ forwards to wrapIOToken(copyFile(src, dst, _)); }

abstract production touchFileM
top::IOMonad<Unit> ::= file::String
{ forwards to wrapIOToken(touchFile(file, _)); }
