grammar test:lexer_b;

lexer class B;