grammar silver:host:env;

-- concrete syntax
exports silver:definition:env:parser;
exports silver:definition:core:env_parser;
exports silver:definition:concrete_syntax:env_parser;

-- symbols
exports silver:definition:env;

