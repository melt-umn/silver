grammar silver:analysis;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Analysis\nmenu_title: Analysis\nmenu_weight: 100\n---"
@}

