grammar simple:host ;

exports simple:terminals ;
exports simple:concretesyntax ;
exports simple:abstractsyntax ;

import simple:concretesyntax only Root_c ;

