grammar silver:compiler:extension:list;

imports silver:compiler:definition:type;
imports silver:compiler:definition:env;
imports silver:compiler:definition:core;

exports silver:compiler:extension:list:java with silver:compiler:translation:java:type;


