grammar silver:compiler:translation:java;

exports silver:compiler:translation:java:core;
exports silver:compiler:translation:java:type;

exports silver:compiler:translation:java:driver;

