grammar silver:extension:monad;

imports silver:definition:core;
imports silver:definition:type:syntax;

imports silver:definition:env;
imports silver:definition:type;

imports silver:extension:convenience;
imports silver:modification:lambda_fn;
imports silver:modification:let_fix;

--import silver:util;