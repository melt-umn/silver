@@{-
    @config grammarWeight -10-}
@{-
  - 
  - Docs for B/bar
  -
  - Second stanza.
  -}
function bar
Integer ::= {return 0;}
