grammar copper_features;

imports silver:testing ;
imports lib:extcore ;

mainTestSuite copper_tests ;

{- Needed: 
layout tests
precedence / associativity tests
lexer classes & dominates submits tests
production precedence / operator tests
-}
