grammar silver:analysis:typechecking:concrete_syntax;

