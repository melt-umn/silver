grammar silver:modification:let_fix;

attribute defaultInheritedAnnos occurs on AssignExpr;