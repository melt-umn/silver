grammar silver:compiler:extension:datalog;

imports silver:core;
imports silver:compiler:analysis:typechecking:core;
imports silver:compiler:definition:core;
imports silver:compiler:definition:env;
imports silver:compiler:definition:type;
imports silver:compiler:definition:type:syntax;
imports silver:compiler:extension:patternmatching;
imports silver:compiler:extension:silverconstruction;
imports silver:compiler:modification:defaultattr;
