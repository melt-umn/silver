grammar copper_features:mdatests;

import copper_features:mdatests:host;
import copper_features:mdatests:ext;

copper_mda test(doParse) {
  copper_features:mdatests:ext;
}


