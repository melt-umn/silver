grammar silver_features:cond:a;

exports silver_features:cond:c with silver_features:cond:b;
