grammar implicit_monads;

imports silver:testing;

mainTestSuite implicit_monad_tests;

{-
  I'm putting this in its own test suite beacuse including it in
  silver_features was causing the testing to stack overflow.
-}

