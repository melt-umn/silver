grammar silver:compiler:extension:patternmatching;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Pattern Matching\nmenu_title: Pattern Matching\nmenu_weight: 100\n---"
@}
