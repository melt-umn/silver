grammar silver:compiler:modification;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Modification\nmenu_title: Modification\nmenu_weight: 100\n---"
@}

