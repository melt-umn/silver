grammar silver_features ;

imports silver:testing ;
imports lib:extcore ;

import silver_features:defs ;

mainTestSuite silver_tests ;

