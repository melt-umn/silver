grammar silver:extension:doc:core;

imports silver:definition:core;
imports silver:definition:type:syntax;

imports silver:definition:env;
imports silver:definition:type;

imports silver:extension:convenience;

import silver:util;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Core\nmenu_title: Core\nmenu_weight: 100\n---"
@}
