grammar silver:analysis:typechecking:driver;
export silver:analysis:typechecking:driver;