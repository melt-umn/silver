grammar silver:modification:impide;

imports silver:definition:core;
imports silver:definition:env;

imports silver:definition:concrete_syntax;
imports silver:modification:copper;

imports silver:definition:concrete_syntax:ast;
imports silver:modification:impide:cstast;

imports ide;
