grammar silver:compiler:definition:concrete_syntax:copper;

-- edu.umn.cs.melt.copper.compiletime.spec.grammarbeans.GrammarElement
type GrammarElement foreign;

-- edu.umn.cs.melt.copper.compiletime.spec.grammarbeans.DisambiguationFunction

-- edu.umn.cs.melt.copper.compiletime.spec.grammarbeans.GrammarSymbol

-- edu.umn.cs.melt.copper.compiletime.spec.grammarbeans.OperatorClass

-- edu.umn.cs.melt.copper.compiletime.spec.grammarbeans.ParserAttribute

-- edu.umn.cs.melt.copper.compiletime.spec.grammarbeans.Production

-- edu.umn.cs.melt.copper.compiletime.spec.grammarbeans.TerminalClass
