@@{-Doc foo foo-}

@{--}
function foo
Integer ::=
{ return 0; }

function undocumented
Integer ::=
{ return 0; }

