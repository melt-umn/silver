grammar tutorials:dc ;

-- Concrete Syntax --
---------------------

