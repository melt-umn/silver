grammar xrobots:terminals ;

-- type keywords

terminal Int_t 'int' dominates { Id_t } ;
terminal Boolean_t  'boolean'  dominates { Id_t } ;
terminal Real_t  'real' dominates { Id_t } ;
terminal Float_t  'float' dominates { Id_t };
terminal String_t  'string' dominates { Id_t };

