imports doctest:nonsplit:childsplit:anotherlevel;

@@{-Doc in X.sv-}

@@{-Second doc in X.sv-}
@@{-@config title "File X"-}