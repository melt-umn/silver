grammar tutorials:xrobots:host ;

--exports tutorials:xrobots:terminals ;
--exports tutorials:xrobots:concretesyntax ;
--exports tutorials:xrobots:abstractsyntax ;

import tutorials:xrobots:concretesyntax only Root_c ;

