
-- The point of this file is to ensure comments are parsed properly.

equalityTest(ca,1,Integer,silver_tests);
equalityTest(cb,1,Integer,silver_tests);
equalityTest(cc,1,Integer,silver_tests);
equalityTest(cd,1,Integer,silver_tests);
equalityTest(ce,1,Integer,silver_tests);
equalityTest(cf,1,Integer,silver_tests);
equalityTest(cg,1,Integer,silver_tests);
equalityTest(ch,1,Integer,silver_tests);
equalityTest(ci,1,Integer,silver_tests);
equalityTest(cj,1,Integer,silver_tests);


{- testing -}

global ca::Integer = 1;

-- testing

global cb::Integer = 1;

{- testing
-}

global cc::Integer = 1;

{- -- -}
global cd::Integer = 1;

{--}
global ce::Integer = 1;

{---}
global cf::Integer = 1;

{----}

global cg::Integer = 1;

{-


testibn


-}

global ch::Integer = 1;

{-
 -
 - hi
 -}
 
global ci::Integer = 1;

 
{-{--}

global cj::Integer = 1;


