grammar lib:lsp;

exports lib:lsp:codeAction;
exports lib:lsp:codeLens;
exports lib:lsp:color;
exports lib:lsp:completion;
exports lib:lsp:constants;
exports lib:lsp:diagnostic;
exports lib:lsp:document;
exports lib:lsp:document:highlight;
exports lib:lsp:document:link;
exports lib:lsp:document:synchronization;
exports lib:lsp:executeCommand;
exports lib:lsp:files;
exports lib:lsp:folding;
exports lib:lsp:formatting;
exports lib:lsp:hover;
exports lib:lsp:goTo;
exports lib:lsp:initialization;
exports lib:lsp:json;
exports lib:lsp:messages;
exports lib:lsp:references;
exports lib:lsp:registration;
exports lib:lsp:rename;
exports lib:lsp:shutdown;
exports lib:lsp:signatureHelp;
exports lib:lsp:symbols;
exports lib:lsp:workspace;
