grammar lib:stringmap;

{@config
  no-doc:"true"
@}

