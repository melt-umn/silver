grammar tutorials:expr:terminals ;

terminal Int_t 'int' dominates { Id_t } ;
terminal Boolean_t  'boolean'  dominates { Id_t } ;

