grammar lib:extcore;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Extended Core\nmenu_title: Extended Core\nmenu_weight: 100\n---"
@}

