
imports lib:lsp:json;
imports lib:lsp:document;
imports lib:lsp;
