grammar lib:monto;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Monto\nmenu_title: Monto\nmenu_weight: 100\n---"
@}

