
terminal Single_t 'single';


equalityTest( 'single'.lexeme, "single", String, silver_tests );
