grammar silver:modification:copper;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Copper\nmenu_title: Copper\nmenu_weight: 100\n---"
@}

