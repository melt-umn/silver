grammar silver:translation:java:type:io;
export silver:translation:java:type:io;


