grammar silver:compiler:extension:scopegraphs;

imports silver:compiler:definition:core;
imports silver:compiler:definition:type;

--imports silver:regex:concrete_syntax;
--imports silver:regex as abs;