grammar silver:modification:let_fix;

build silver:modification:let_fix:java with silver:translation:java;

