grammar xrobots:host ;

--exports tutorials:xrobots:terminals ;
--exports tutorials:xrobots:concretesyntax ;
--exports tutorials:xrobots:abstractsyntax ;

import xrobots:concretesyntax only Root_c ;

