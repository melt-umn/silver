
imports lib:lsp;
