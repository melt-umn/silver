@@{-

@config excludeFile

Docs in A.sv-}