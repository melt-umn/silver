grammar silver:definition:type:syntax;


terminal Boolean_tkwd    'Boolean'   lexer classes {TYPE,RESERVED};
terminal Decorated_tkwd  'Decorated' lexer classes {TYPE,RESERVED};
terminal Float_tkwd      'Float'     lexer classes {TYPE,RESERVED};
terminal Integer_tkwd    'Integer'   lexer classes {TYPE,RESERVED};
terminal String_tkwd     'String'    lexer classes {TYPE,RESERVED};


