grammar silver:extension:ideinterface;

imports silver:definition:env;
imports silver:definition:core;
imports silver:definition:type;
imports silver:definition:regex;
imports silver:definition:concrete_syntax;
imports silver:definition:concrete_syntax:ast;

nonterminal IdeInterfaceRoot;
