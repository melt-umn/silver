grammar core:reflect;

function reflect
AST ::= x::a
{
  return error("Foreign function");
} foreign {
  "java" : return "(common.Reflection.reflect(%x%))";
}

function reflectTypeName
Maybe<String> ::= x::a
{
  return error("Foreign function");
}{- foreign {
  "java" : return "(common.Reflection.reflectTypeName(%x%))";
}-}
