grammar silver:compiler:modification:autocopyattr;

imports silver:compiler:definition:env;
imports silver:compiler:definition:core;
imports silver:compiler:definition:type;
imports silver:compiler:definition:type:syntax;

exports silver:compiler:modification:autocopyattr:java with silver:compiler:translation:java:core;
exports silver:compiler:modification:autocopyattr:convenience with silver:compiler:extension:convenience;

