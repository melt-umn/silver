grammar simple:extensions:matrix;

imports lib:lang;
imports simple:concretesyntax as cst;
imports simple:abstractsyntax;


terminal Matrix 'Matrix' lexer classes { KEYWORDS };
terminal LBrack '[';
terminal RBrack ']';


