grammar silver:extension:list;

