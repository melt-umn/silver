function sub
Integer ::= a::Integer b::Integer
{
	return add(a, -b);
}