grammar tutorials:simple:host ;

exports tutorials:simple:terminals ;
exports tutorials:simple:concretesyntax ;
exports tutorials:simple:abstractsyntax ;

import tutorials:simple:concretesyntax only Root_c ;

