grammar silver:compiler:extension:easyterminal;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Easy Terminal\nmenu_title: Easy Terminal\nmenu_weight: 100\n---"
@}

