grammar silver:xml:ast;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Abstract Syntax Tree\nmenu_title: AST\nmenu_weight: 100\n---"
@}

