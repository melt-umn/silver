grammar tutorials:simple:abstractsyntax ;

nonterminal Root ;
