grammar lib:lsp:hover;

imports lib:lsp;
