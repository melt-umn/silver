
imports lib:lsp;
--imports lib:lsp:json;
--imports lib:lsp:document;
--imports lib:lsp:diagnostic;
--imports lib:lsp:executeCommand;
--imports lib:lsp:workspace;
