grammar silver:modification:collection;

imports silver:definition:env;
imports silver:definition:core;
imports silver:definition:type;

exports silver:modification:collection:java with silver:translation:java:core;

