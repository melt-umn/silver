grammar silver:analysis:typechecking:command;
export silver:analysis:typechecking:command;
