grammar silver:definition:core;

{--
 - The grammar containing this tree.
 -}
autocopy attribute grammarName :: String;
