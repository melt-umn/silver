grammar silver:compiler:modification:copper_mda;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Copper MDA\nmenu_title: Copper MDA\nmenu_weight: 100\n---"
@}

