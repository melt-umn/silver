grammar silver:compiler:extension:abella_compilation:abella;

imports silver:compiler:definition:core;
imports silver:compiler:definition:env;
imports silver:compiler:definition:type;

