grammar silver:modification:ffi;

exports silver:modification:ffi:java with silver:translation:java;

