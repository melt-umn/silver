grammar silver:xml;

{@config
  header:"---\nlayout: sv_wiki\ntitle: XML\nmenu_title: XML\nmenu_weight: 100\n---"
@}

