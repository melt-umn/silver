grammar core;

nonterminal UnitT;

abstract production unit
top::UnitT ::=
{}