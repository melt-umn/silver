grammar silver:extension:bidirtransform;

synthesized attribute rewriteRules::[Decorated RewriteRule];
synthesized attribute outputStmt::(Expr ::= Expr);
synthesized attribute restoreStmt::(Expr ::= Expr);
synthesized attribute inputType::Type;
synthesized attribute inputProduction::RewriteProduction;
synthesized attribute hasProduction::Boolean;
synthesized attribute shouldRestore::Boolean;
synthesized attribute decSig::Decorated NamedSignature;
synthesized attribute rhsType::Maybe<TypeExpr>;

nonterminal RewriteRuleList with rewriteRules, env, errors, location, absGroup, cncGroup, pp, downSubst, upSubst, finalSubst, config;
nonterminal RewriteRule with inputType, inputProduction, hasProduction, typerep, outputStmt, restoreStmt, shouldRestore, env, errors, location, absGroup, cncGroup, pp, downSubst, upSubst, finalSubst, config;
nonterminal RewriteProduction with name, inputNames, typerep, env, errors, location, absGroup, cncGroup, pp, config, decSig;
nonterminal RewriteProductionArgs with inputNames, errors, pp, config;
nonterminal RewriteArrow with shouldRestore, rhsType;
nonterminal OptRHSType with rhsType;

terminal RestoreArrow_t '~~>' lexer classes {SPECOP};

concrete production rewriteRuleCons
rrl::RewriteRuleList ::= Vbar_kwd l::RewriteRule r::RewriteRuleList
{
    l.downSubst = rrl.downSubst;
    r.downSubst = l.upSubst;
    rrl.upSubst = r.upSubst;
    l.finalSubst = r.upSubst;
    r.finalSubst = l.finalSubst;

    rrl.pp = "| " ++ l.pp ++ r.pp;

    rrl.errors := l.errors ++ r.errors;
    rrl.rewriteRules = r.rewriteRules ++ [l];
    
    -- error check: is the exact rule l found in r?
    -- equality checking is non trivial so we aren't doing this
    -- rrl.errors <- if !containsBy(\ a::RewriteRule b::RewriteRule -> eq(a,b), l, r.rewriteRules) then []
    --               else [err(rrl.location, "Duplicate rewrite rule definition")];

}

concrete production rewriteRuleSingle
rrl::RewriteRuleList ::= Vbar_kwd rule::RewriteRule 
{
    rule.downSubst = rrl.downSubst;
    rrl.upSubst = rule.upSubst;
    rule.finalSubst = rrl.upSubst;

    rrl.pp = "| " ++ rule.pp;

    rrl.rewriteRules = [rule];
    rrl.errors := rule.errors;
}

-- rewrite a production as another production,
-- recursing on restored elements
concrete production rewriteRuleProd
rule::RewriteRule ::= prd::RewriteProduction arr::RewriteArrow e::Expr
{
    rule.pp = prd.pp ++ "~~>" ++ e.pp;

    e.downSubst = rule.downSubst;
    rule.upSubst = e.upSubst;
    e.finalSubst = rule.upSubst;
    e.defaultInheritedAnnos = [];

    local rhsType::Type = case arr.rhsType of 
        | just(t) -> t.typerep
        | nothing() -> e.typerep
    end;      

    forwards to rewriteRule(e, "", prd.typerep, rhsType, 
        prd, true, arr.shouldRestore, location=rule.location);
}

-- rewrite a  type as another type through plugging it into
-- an expression
concrete production rewriteRuleType
rule::RewriteRule ::= name::QName '::' t::TypeExpr arr::RewriteArrow  e::Expr
{
    rule.pp = name.pp ++ "::" ++ t.pp ++ "~~>" ++ e.pp;

    -- I shouldn't need to have to redefine this, as the forward defines this, but I do.
    e.downSubst = rule.downSubst;
    rule.upSubst = e.upSubst;
    e.finalSubst = rule.upSubst;
    e.defaultInheritedAnnos = [];     

    local rhsType::Type = case arr.rhsType of 
        | just(t) -> t.typerep
        | nothing() -> e.typerep
    end;
    
    forwards to rewriteRule(e, name.name, t.typerep, rhsType, 
      emptyRewriteProduction(location=rule.location), false, arr.shouldRestore, location=rule.location);
}

concrete production shortRewriteArrow
arr::RewriteArrow ::= '->' opt::OptRHSType 
{
    arr.shouldRestore = false;
    arr.rhsType = opt.rhsType;
}

concrete production longRewriteArrow
arr::RewriteArrow ::= '~~>' opt::OptRHSType 
{
    arr.shouldRestore = true;
    arr.rhsType = opt.rhsType;
}

concrete production oneRHSType
opt::OptRHSType ::= Vbar_kwd t::TypeExpr Vbar_kwd
{
    opt.rhsType = just(t);
}

concrete production noRHSType
opt::OptRHSType ::= 
{
    opt.rhsType = nothing();
}

abstract production rewriteRule
rule::RewriteRule ::= rhs::Expr inName::String inType::Type outType::Type inProd::RewriteProduction hasProd::Boolean restore::Boolean
{
    rhs.downSubst = rule.downSubst;
    rule.upSubst = rhs.upSubst;
    rhs.finalSubst = rule.upSubst;

    rhs.defaultInheritedAnnos = [];

    rule.errors := []; -- We explicitly ignore rhs errors here
    rule.errors <- inProd.errors;
    -- rule.errors <- [err(rule.location, "rwRule:" ++ rhs.pp ++ "in,out: " ++ inType.typeName ++ ", " ++ outType.typeName)];

    local rhsNs::Maybe<Decorated NamedSignature> = case rhs of 
        | application(e,_,_,_,_,_) -> case e of
            | baseExpr(qn) -> just(head(getProdFromGroups(qn.name, rule.absGroup, rule.cncGroup)))
            | _ -> nothing()
        end
        | _ -> nothing()
    end;

    rule.hasProduction = hasProd;
    rule.typerep = outType;
    rule.inputType = inType;
    rule.inputProduction = inProd;
    rule.shouldRestore = restore;
    rule.outputStmt = if !hasProd
        then (\ e::Expr -> 
            fillExpr(rhs, [e], [inName], location=e.location))
        else (\ e::Expr ->
            case e of application(_, _, aexpr, _, _, _) -> 
                fillExpr(rhs, pullOutAppExprs(aexpr, top.env), inProd.inputNames, location=e.location)
            end
        );

    rule.restoreStmt = (\ e::Expr ->
            case e of application(_, _, aexpr, _, _, _) -> 
                restoreExpr(rhs, pullOutAppExprs(aexpr, top.env), inProd.inputNames, rhsNs.fromJust, location=e.location)
            end
        );
}