grammar test:term_b;

terminal B_t 'AA';