grammar silver:compiler:extension:deriving;

imports silver:compiler:definition:core;
imports silver:compiler:definition:env;
imports silver:compiler:definition:type;
imports silver:compiler:definition:type:syntax;
imports silver:compiler:modification:collection;
imports silver:compiler:modification:lambda_fn;
imports silver:compiler:modification:primitivepattern;
imports silver:compiler:metatranslation;
