grammar silver:modification:autocopyattr;

imports silver:definition:env;
imports silver:definition:core;
imports silver:definition:type;
imports silver:definition:type:syntax;

exports silver:modification:autocopyattr:java with silver:translation:java:core;
exports silver:modification:autocopyattr:convenience with silver:extension:convenience;

