@@{-Doc in Y.sv-}
@@{-@config split
    @config title "File Y"-}