grammar silver:compiler:extension:implicit_monads;
