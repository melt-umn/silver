grammar silver:compiler:definition;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Definition\nmenu_title: Definition\nmenu_weight: 100\n---"
@}

