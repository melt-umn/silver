grammar silver:compiler:extension:abella_compilation:encoding;

--imports silver:compiler:definition:env;
--imports silver:compiler:definition:core;

imports silver:compiler:definition:core;
imports silver:compiler:definition:type;
imports silver:compiler:definition:type:syntax;
imports silver:compiler:extension:list;

imports silver:compiler:definition:concrete_syntax;
imports silver:compiler:modification:ffi;
imports silver:compiler:extension:autoattr;
imports silver:compiler:modification:defaultattr;
imports silver:compiler:modification:copper;
imports silver:compiler:modification:copper_mda;
imports silver:compiler:definition:flow:syntax;
imports silver:compiler:modification:collection;
imports silver:compiler:definition:env;

imports silver:compiler:extension:abella_compilation:abella;

