grammar lib:errors;

{@config
  no-doc:"true"
@}

