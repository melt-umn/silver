grammar recTy;

exports host;

type RecErr = RecErr;

parser extendedParser :: Root {
    host;
    recTy;
} 