grammar silver_features:cond:b;

-- empty, dummy grammar.
