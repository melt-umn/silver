grammar silver:compiler:extension:doc;

exports silver:compiler:extension:doc:core;
exports silver:compiler:extension:doc:driver;



