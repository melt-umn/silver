grammar silver:translation:java:concrete_syntax;

