grammar silver:util;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Utilities\nmenu_title: Util\nmenu_weight: 100\n---"
@}

