grammar silver:extension;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Extensions\nmenu_title: Extensions\nmenu_weight: 100\n---"
@}

