grammar silver:modification:let_fix;

imports silver:definition:core;
imports silver:definition:env;
imports silver:definition:type;
imports silver:definition:type:syntax;
imports silver:analysis:typechecking;
imports silver:analysis:typechecking:core;

exports silver:modification:let_fix:java with silver:translation:java;

