@@{-

@config excludeFile

Docs in Excluded.sv-}