@@{-Docs in Second.sv-}