grammar silver:core;

equality attribute isEqualTo, isEqual;
