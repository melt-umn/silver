grammar silver_features:cond:c;

exports silver_features:cond:d;

global aVal :: Integer = 1;

