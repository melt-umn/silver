grammar silver:extension:implicit_monads;

imports silver:definition:core;
imports silver:definition:type:syntax;
imports silver:definition:flow:driver;
imports silver:definition:flow:ast;
imports silver:driver:util;

imports silver:definition:env;
imports silver:definition:type;

imports silver:extension:convenience;
imports silver:extension:patternmatching;

imports silver:modification:lambda_fn;
imports silver:modification:let_fix;
