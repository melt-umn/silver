
nonterminal Bar;

synthesized attribute bs :: String occurs on Bar;
inherited attribute bi :: String occurs on Bar;

abstract production barBar
t::Bar ::= {}


