@@{-Doc foo foo-}

@{-Docs on foo-}
function foo
Integer ::=
{ return 0; }

function undocumented
Integer ::=
{ return 0; }

function undocumented2
Integer ::=
{ return 0; }

