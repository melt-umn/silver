
terminal Propagate_kwd 'propagate' lexer classes {KEYWORD,RESERVED};
terminal Functor_kwd   'functor' lexer classes {KEYWORD,RESERVED};
terminal Monoid_kwd    'monoid' lexer classes {KEYWORD,RESERVED};
