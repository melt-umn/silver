grammar tutorials:hello;

function main 
IOVal<Integer> ::= largs::[String] ioin::IO
{
  return ioval(print(" World!\n",
                 print("Hello", ioin)),
               0);
}
