grammar core;

exports core:monad;