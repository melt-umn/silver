imports doctest:nonsplit:childsplit;

@{-
  - Docs for A/foo
  -}
function foo
Integer ::= {return 0;}