grammar silver:modification:impide:spec;

imports silver:definition:core;
imports silver:definition:env;

imports silver:definition:concrete_syntax;
imports silver:modification:copper;

imports silver:definition:concrete_syntax:ast;
imports silver:modification:impide:cstast;
imports silver:modification:impide;

imports silver:translation:java:core only makeClassName, makeParserName;

