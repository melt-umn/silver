grammar monto:concretesyntax;

imports monto:abstractsyntax as abs;

-- Used to build the abstract syntax tree from the concrete syntax tree
synthesized attribute ast<a>::a;
