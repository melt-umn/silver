package test:prod_b;

exports test:nonterm_b;

concrete production B_p
B ::=
{    
}