imports lib:lsp;
