grammar silver:modification:typedecl;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Type Declarations\nmenu_title: Type Declarations\nmenu_weight: 100\n---"
@}

