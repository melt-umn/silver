grammar silver:translation:java:type:anytype;
export silver:translation:java:type:anytype;
