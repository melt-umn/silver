grammar silver:compiler:modification:let_fix;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Let Fix\nmenu_title: Let Fix\nmenu_weight: 100\n---"
@}

