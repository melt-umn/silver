grammar lib:lsp:workspace;

imports lib:lsp:document;
imports lib:lsp:json;
imports lib:lsp;
imports lib:lsp:symbols;
