grammar silver:extension:templating:syntax;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Syntax\nmenu_title: Syntax\nmenu_weight: 100\n---"
@}

