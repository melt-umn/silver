grammar silver:definition:core;

import silver:definition:env;

concrete production qNameId
top::QName ::= id::Name
{
  top.name = id.name;
  top.pp = id.pp;
  top.location = id.location;
  
  top.lookupValue = decorate customLookup("value", getValueDcl, top) with { env = top.env; };
  top.lookupType = decorate customLookup("type", getTypeDcl, top) with { env = top.env; };
  top.lookupAttribute = decorate customLookup("attribute", getAttrDcl, top) with { env = top.env; };
}

concrete production qNameCons
top::QName ::= id::Name ':' qn::QName
{
  top.name = id.name ++ ":" ++ qn.name;
  top.pp = id.pp ++ ":" ++ qn.pp;
  top.location = loc(top.file, $2.line, $2.column);
  
  top.lookupValue = decorate customLookup("value", getValueDcl, top) with { env = top.env; };
  top.lookupType = decorate customLookup("type", getTypeDcl, top) with { env = top.env; };
  top.lookupAttribute = decorate customLookup("attribute", getAttrDcl, top) with { env = top.env; };
}

synthesized attribute lookupValue :: Decorated QNameLookup occurs on QName;
synthesized attribute lookupType :: Decorated QNameLookup occurs on QName;
synthesized attribute lookupAttribute :: Decorated QNameLookup occurs on QName;

nonterminal QNameLookup with fullName, typerep, errors, env, dcls, dcl;

abstract production customLookup
top::QNameLookup ::= lookupName::String lookupFunc::Function([Decorated DclInfo] ::= String Decorated Env) q::Decorated QName 
{
  top.dcls = lookupFunc(q.name, top.env);
  top.dcl = head(top.dcls);
  
  top.fullName = top.dcl.fullName;
  
  top.typerep = if null(top.dcls)
                then topTypeRep()
                else head(top.dcls).typerep;
  
  top.errors := (if null(top.dcls)
                  then [err(q.location, "Undeclared " ++ lookupName ++ " '" ++ q.name ++ "'.")]
                  else [])
             ++ (if length(top.dcls) > 1
                  then [err(q.location, "Ambiguous reference to " ++ lookupName ++ " '" ++ q.name ++ "'. Possibilities are:\n" ++ printPossibilities(top.dcls))] 
                  else []);
}

function printPossibilities
String ::= lst::[Decorated DclInfo]
{
  local attribute dcl :: Decorated DclInfo;
  dcl = head(lst);
  
  -- TODO: perhaps some way of including types, when they are relevant (attributes, values)
  return if null(lst) then ""
         else ("\t" ++ dcl.fullName ++ " (" ++ dcl.sourceLocation.fileName ++ ":" ++ toString(dcl.sourceLocation.line) ++ ")\n")
              ++ printPossibilities(tail(lst));
}

