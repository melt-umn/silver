grammar silver:modification:autocopyattr;

exports silver:modification:autocopyattr:java with silver:translation:java:core;
exports silver:modification:autocopyattr:convenience with silver:extension:convenience;

