grammar silver:extension:list;

imports silver:definition:type;
imports silver:definition:env;
imports silver:definition:core;

exports silver:extension:list:java with silver:translation:java:type;

