grammar silver_features:cond:a;

build silver_features:cond:c with silver_features:cond:b;
