grammar silver:compiler:extension:doc:core;

imports silver:compiler:definition:core;
imports silver:compiler:definition:type:syntax;

imports silver:compiler:definition:env;
imports silver:compiler:definition:type;

imports silver:compiler:extension:convenience hiding ProdVBar;

imports silver:util:treemap as tm;
