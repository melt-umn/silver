grammar silver:extension:list;

build silver:extension:list:java with silver:translation:java;

