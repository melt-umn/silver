grammar lib:lsp:document;

imports lib:lsp;
