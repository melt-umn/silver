grammar silver_features:cond:c;

global aVal :: Integer = 1;

