
imports lib:lsp;
imports lib:lsp:json;
imports lib:lsp:document;
imports core hiding Location;
