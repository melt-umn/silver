grammar silver:definition;
export silver:definition;

