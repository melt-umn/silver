grammar silver:modification:collection;

build silver:modification:collection:java with silver:translation:java;

