grammar silver:analysis:binding:driver;
export silver:analysis:binding:driver;