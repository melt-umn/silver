grammar silver:extension:list;

exports silver:extension:list:java with silver:translation:java;

