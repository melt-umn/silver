grammar stdlib:rewrite;

exports stdlib:rewrite:expreval;
