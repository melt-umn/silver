
type DocumentSelector = [DocumentFilter];
