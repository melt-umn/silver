grammar silver:extension:doc:core;

nonterminal DocItem;

abstract production commentDocItem
top::DocItem ::= c::CommentItem
{}


