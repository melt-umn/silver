@@{-Docs in Second.sv-}

function exFn
Boolean ::= {return true;}