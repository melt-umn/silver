grammar silver:compiler:extension:datalog;
