@@{-Doc foo foo-}

@{--}
function foo
Integer ::=
{ return 0; }