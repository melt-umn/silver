-- This will be used in issue #17.
-- The following generates an inappropriate error message.
-- The intTestProd is defined in FuncProdTypes.sv
-- equalityTest ( intTestProd(0), 0, Integer, silver_tests ) ;
