grammar lib:system;

{@config
  header:"---\nlayout: sv_wiki\ntitle: System\nmenu_title: System\nmenu_weight: 100\n---"
@}

