grammar silver:core;

data nonterminal Unit;

abstract production unit
top::Unit ::=
{}