grammar silver:analysis:typechecking:type:anytype;
export silver:analysis:typechecking:type:anytype;
