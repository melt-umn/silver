grammar silver:compiler:composed;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Composed\nmenu_title: Composed\nmenu_weight: 100\n---"
@}

