grammar tutorials:dc ;
