grammar lib:lsp:json;

parser jsonParser :: JSONText {
  lib:lsp:json;
} 
