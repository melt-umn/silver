grammar silver:modification:annotation;


