grammar silver:modification:collection:java;
export silver:modification:collection:java;
