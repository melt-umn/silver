imports lib:lsp;
imports lib:lsp:codeAction;
imports lib:lsp:codeLens;
imports lib:lsp:completion;
imports lib:lsp:constants;
imports lib:lsp:document;
imports lib:lsp:document:link;
imports lib:lsp:executeCommand;
imports lib:lsp:formatting;
imports lib:lsp:json;
imports lib:lsp:rename;
imports lib:lsp:signatureHelp;
imports lib:lsp:workspace;
