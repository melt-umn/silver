@@{-Content-}