grammar silver:modification:origintracking;

imports silver:definition:type;
imports silver:definition:type:syntax;
imports silver:definition:env;
imports silver:definition:core;

imports silver:translation:java:core;
imports silver:translation:java:type;

-- imports silver:extension:otx:childruntime; -- So we can make sure it builds