imports silver:reflect;