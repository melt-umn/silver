grammar silver:analysis:binding:command;
export silver:analysis:binding:command;