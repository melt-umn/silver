
imports lib:lsp:json;
imports lib:lsp;
imports lib:lsp:document;
