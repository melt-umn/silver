
imports lib:lsp;
imports core hiding Location;
