grammar core;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Core\nmenu_title: Core library\nmenu_weight: 20\n---"

  split-files: true
@}

