grammar core:monad;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Monad support\nmenu_title: Monads\nmenu_weight: 50\n---"
@}
