grammar silver:extension:functorattrib;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Functor Attributes\nmenu_title: Functor Attributes\nmenu_weight: 100\n---"
@}

