grammar silver:compiler:modification:autocopyattr;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Autocopy Attribute\nmenu_title: Autocopy Attribute\nmenu_weight: 100\n---"
@}
