grammar silver:extension:list;

imports silver:definition:type;
imports silver:definition:env;
imports silver:definition:core;

exports silver:extension:list:java with silver:translation:java:type;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Lists\nmenu_title: Lists\nmenu_weight: 100\n---"
@}
