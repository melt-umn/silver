grammar silver:extension:autoattr;

terminal Propagate_kwd 'propagate' lexer classes {KEYWORD,RESERVED};
terminal Excluding_kwd 'excluding' lexer classes {KEYWORD};
terminal Thread_kwd    'thread'    lexer classes {KEYWORD,RESERVED};

terminal Functor_kwd     'functor'     lexer classes {KEYWORD,RESERVED};
terminal Monoid_kwd      'monoid'      lexer classes {KEYWORD,RESERVED};
terminal Equality_kwd    'equality'    lexer classes {KEYWORD,RESERVED};
terminal Unification_kwd 'unification' lexer classes {KEYWORD,RESERVED};
terminal Threaded_kwd    'threaded'    lexer classes {KEYWORD,RESERVED};
