grammar silver:analysis:typechecking:core;

aspect production defaultClassBodyItem
top::ClassBodyItem ::= id::Name '::' ty::TypeExpr '=' e::Expr ';'
{
  top.errors <-
    if ty.typerep.kindArity > 0
    then [err(ty.location, s"Type ${ty.unparse} is not fully applied, it has kind arity ${toString(ty.typerep.kindArity)}")]
    else [];

  local errCheck1::TypeCheck = check(ty.typerep, e.typerep);
  top.errors <-
    if errCheck1.typeerror
    then [err(e.location, s"Member ${id.name} has expected type ${errCheck1.leftpp}, but the expression has actual type ${errCheck1.rightpp}")]
    else [];
  
  e.downSubst = emptySubst();
  errCheck1.downSubst = e.upSubst;
  e.finalSubst = e.upSubst;
  errCheck1.finalSubst = e.finalSubst;
}
