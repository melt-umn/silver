
grammar monto:abstractsyntax;

{- This file holds attribute declarations for abstract syntax. -}

synthesized attribute value::Integer;
synthesized attribute errors::[String];
synthesized attribute tostring::String;
