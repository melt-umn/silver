grammar lib:system ;

exports lib:system:filenames ;
exports lib:system:ioaction ;
