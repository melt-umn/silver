grammar tutorials:hello;


function main
IO ::= args::String ioin::IO
{
  return print(" World!\n",
           print("Hello", ioin));
}
