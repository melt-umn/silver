grammar silver:modification:impide;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Imp IDE\nmenu_title: Imp IDE\nmenu_weight: 100\n---"
@}

