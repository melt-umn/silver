grammar silver:translation:java;

exports silver:translation:java:core;
exports silver:translation:java:env;
exports silver:translation:java:concrete_syntax;
exports silver:translation:java:type:io;
exports silver:translation:java:type:anytype;

exports silver:translation:java:driver;

