grammar silver:compiler:modification:defaultattr;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Default Attribute\nmenu_title: Default Attribute\nmenu_weight: 100\n---"
@}

