grammar silver:testing;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Testing\nmenu_title: Testing\nmenu_weight: 100\n---"
@}

