import silver:json;

synthesized attribute json :: Json;
