grammar silver:compiler:langserver;

-- This grammar contains helper functions and attributes used in the Silver LSP implementation.
-- For simplicitly, this grammar is imported in the build of the normal compiler for now.

imports silver:compiler:host;
imports silver:compiler:definition:env;

imports silver:util:treemap as map;
