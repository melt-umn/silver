grammar silver:modification:collection;

