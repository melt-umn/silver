grammar silver:compiler:extension:implicit_monads;

imports silver:compiler:definition:core;
imports silver:compiler:definition:type:syntax hiding Unique_t;
imports silver:compiler:definition:flow:driver;
imports silver:compiler:definition:flow:ast;
imports silver:compiler:definition:flow:env;
imports silver:compiler:driver:util;

imports silver:compiler:definition:env;
imports silver:compiler:definition:type;
imports silver:compiler:analysis:typechecking:core;

imports silver:util:cmdargs;

imports silver:compiler:extension:convenience;
imports silver:compiler:extension:patternmatching;
imports silver:compiler:modification:list;

imports silver:compiler:modification:lambda_fn;
imports silver:compiler:modification:let_fix;
imports silver:compiler:modification:primitivepattern;
imports silver:compiler:modification:copper;
