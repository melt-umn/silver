grammar silver:compiler:extension:doc:core;

synthesized attribute body :: String;
synthesized attribute file :: String;
nonterminal CommentItem with body, file;
