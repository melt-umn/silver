grammar silver:modification:primitivepattern;

attribute defaultInheritedAnnos occurs on PrimPattern, PrimPatterns;