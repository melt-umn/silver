grammar core;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Core\nmenu_title: Core\nmenu_weight: 100\n---"
  split-files:"true"
@}

