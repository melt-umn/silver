grammar silver:compiler:definition:concrete_syntax;

imports silver:langutil:lsp as lsp;

imports silver:compiler:definition:core;
imports silver:compiler:definition:type:syntax;

imports silver:compiler:definition:env;
imports silver:compiler:definition:type;

imports silver:compiler:definition:concrete_syntax:ast;

option silver:compiler:modification:copper;
