grammar silver:compiler:modification:primitivepattern;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Primitive Pattern\nmenu_title: Primitive Pattern\nmenu_weight: 100\n---"
@}

