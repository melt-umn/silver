grammar silver:host;

-- concrete syntax from these grammars
exports silver:definition:core;
exports silver:definition:concrete_syntax;
exports silver:definition:type:io;
exports silver:definition:type:higherorder;
exports silver:definition:type:productiontype;
exports silver:definition:type:decorated;
exports silver:definition:type:anytype;

-- symbols
exports silver:analysis:binding:driver;
exports silver:analysis:typechecking:driver;
exports silver:analysis:typechecking:core;
exports silver:analysis:typechecking:concrete_syntax;
exports silver:analysis:typechecking:type:io;
exports silver:analysis:typechecking:type:anytype;

