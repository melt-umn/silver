grammar silver:util;

-- Just import all the subgrammars here, so we have an easy way to build all of them.
imports silver:util:cmdargs;
imports silver:util:deque;
imports silver:util:graph;
imports silver:util:random;
imports silver:util:subprocess;
imports silver:util:treemap;
imports silver:util:treeset;
imports silver:reflect;
