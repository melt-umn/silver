grammar silver:extension:strategyattr;

imports silver:definition:core;
imports silver:definition:env;
imports silver:definition:type;
imports silver:definition:type:syntax;
imports silver:extension:autoattr;
imports silver:extension:patternmatching;
imports silver:extension:list;
--imports silver:extension:rewriting;
imports silver:modification:let_fix;

exports silver:extension:strategyattr:convenience;
