grammar silver:translation:java:driver;

