grammar silver:extension:autoattr;

imports silver:definition:core;
imports silver:definition:env;
imports silver:definition:type;
imports silver:definition:type:syntax;
imports silver:modification:collection;

exports silver:extension:autoattr:convenience;
