grammar silver:extension:polymorphism;

export silver:extension:polymorphism;
export silver:extension:polymorphism:functions;

syntax silver:extension:polymorphism:functions;