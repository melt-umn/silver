grammar silver:extension:doc;

exports silver:extension:doc:core;
exports silver:extension:doc:driver;

{@config
  no-doc:"true"
@}

