grammar lib:lsp:symbols;

imports lib:lsp:document;
imports lib:lsp:json;
imports lib:lsp;
imports core with Location as CoreLocation;
