grammar silver:translation:java:env;

