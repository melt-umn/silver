
terminal PropagateOld_kwd 'propagate_functor' lexer classes {KEYWORD,RESERVED};
