@@{-Content should be in the grammar file-}