grammar lib:lsp;

imports lib:lsp:codeAction;
imports lib:lsp:codeLens;
imports lib:lsp:color;
imports lib:lsp:completion;
imports lib:lsp:constants;
imports lib:lsp:diagnostic;
imports lib:lsp:document;
imports lib:lsp:document:highlight;
imports lib:lsp:document:link;
imports lib:lsp:document:synchronization;
imports lib:lsp:executeCommand;
imports lib:lsp:files;
imports lib:lsp:folding;
imports lib:lsp:formatting;
imports lib:lsp:hover;
imports lib:lsp:goTo;
imports lib:lsp:initialization;
imports lib:lsp:json;
imports lib:lsp:messages;
imports lib:lsp:references;
imports lib:lsp:registration;
imports lib:lsp:rename;
imports lib:lsp:shutdown;
imports lib:lsp:signatureHelp;
imports lib:lsp:symbols;
imports lib:lsp:workspace;
