grammar silver:modification:autocopyattr;

build silver:modification:autocopyattr:java with silver:translation:java;
build silver:modification:autocopyattr:convenience with silver:extension:convenience;
