grammar simple:extensions:matrix;

imports silver:langutil;
imports silver:langutil:pp;
imports simple:concretesyntax as cst;
imports simple:abstractsyntax;


terminal Matrix 'Matrix' lexer classes { KEYWORDS };
terminal LBrack '[';
terminal RBrack ']';


