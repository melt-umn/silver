grammar silver:compiler:extension:deprecation;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Deprecation\nmenu_title: Deprecation\nmenu_weight: 100\n---"
@}
