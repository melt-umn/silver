grammar recTy;

exports host;

type A = A;

parser extendedParser :: Root {
    host;
    recTy;
} 