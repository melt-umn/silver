grammar recNt;

exports host;

nonterminal B<B>;

parser extendedParser :: Root {
    host;
    recNt;
} 