grammar lib:langproc;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Language Processing\nmenu_title: Language Processing\nmenu_weight: 100\n---"
@}

