grammar silver:analysis:typechecking:core;

