grammar silver:driver;
import silver:definition:core;
import silver:definition:env;
import silver:util;
import silver:util:command;

synthesized attribute code :: Integer;
synthesized attribute order :: Integer;
inherited attribute ioIn :: IO;
synthesized attribute ioOut :: IO;

nonterminal Unit with ioIn, io, code, order;

aspect production run
top::RunUnit ::= iIn::IO args::String
{
  preOps <- [checkSilverHome(silverhome), checkSilverGen(silvergen)];
  preOps <- if a.displayVersion then [printVersion()] else [];
  postOps <- [doInterfaces(depAnalysis.compiledList, silvergen)];
}

function runAll
IOVal<Integer> ::= i::IO l::[Unit]
{
  local attribute now :: Unit;
  now = head(l);
  now.ioIn = i;

  return  if null(l) 
	  then ioval(i, 0)
	  else if now.code != 0
	       then ioval(now.io, now.code)
	       else runAll(now.io, tail(l));
}

abstract production checkSilverHome
top::Unit ::= s::String
{
  local attribute problem :: Boolean;
  problem = s == "/";

  top.io = if problem then print("Missing SILVER_HOME. Installation problem?\n",top.ioIn) else top.ioIn;
  top.code = if problem then 1 else 0;
  top.order = 0;
}

abstract production checkSilverGen
top::Unit ::= s::String
{
  local attribute problem :: Boolean;
  problem = s == "/";

  top.io = if problem then print("Missing SILVER_GEN or -G <path>. A location to store intermediate files is necessary.\n",top.ioIn) else top.ioIn;
  top.code = if problem then 1 else 0;
  top.order = 0;
}

abstract production printVersion
top::Unit ::= 
{
  top.order = 0;
  top.io = print("Silver Version 0.8 pre-release\n", top.ioIn);
  top.code = -1;
}

abstract production doInterfaces
top::Unit ::= u::[Decorated RootSpec] genPath::String
{
  top.order = 3;
  top.io = writeInterfaces(print("Writing updated interface files\n", top.ioIn), u, genPath);
  top.code = 0;
}

function writeInterfaces
IO ::= iIn::IO r::[Decorated RootSpec] genPath::String
{
  return if null(r) then iIn else writeInterfaces(writeInterface(iIn, head(r), genPath), tail(r), genPath);
}

function writeInterface
IO ::= iIn::IO r::Decorated RootSpec genPath::String
{
  local attribute pathName :: String;
  pathName = genPath ++ "src/" ++ substitute("/", ":", r.impliedName) ++ "/";

  local attribute mkio :: IO;
  mkio = mkdir(pathName, iIn).io;
  
  local attribute pr :: IO;
  pr = print("\t[" ++ r.impliedName ++ "]\n", mkio);
  
  local attribute rm :: IO;
  rm = deleteStaleData(pr, genPath, r.impliedName);
  
  local attribute wr :: IO;
  wr = writeFile(pathName ++ "Silver.svi", r.unparse, rm);
  
  return wr;
}

function deleteStaleData
IO ::= iIn::IO genPath::String gram::String
{
  local attribute srcPath :: String;
  srcPath = genPath ++ "src/" ++ substitute("/", ":", gram) ++ "/";

  local attribute binPath :: String;
  binPath = genPath ++ "bin/" ++ substitute("/", ":", gram) ++ "/";
  
  local attribute srcFiles :: IOVal<[String]>;
  srcFiles = listContents(srcPath, iIn);
  
  local attribute binFiles :: IOVal<[String]>;
  binFiles = listContents(binPath, srcFiles.io);
  
  return deleteStaleDataFiles( deleteStaleDataFiles( binFiles.io, binPath, binFiles.iovalue), srcPath, srcFiles.iovalue);
         
}
function deleteStaleDataFiles
IO ::= iIn::IO path::String files::[String]
{
  local attribute isf :: IOVal<Boolean>;
  isf = isFile(path ++ head(files), iIn);
  
  return if null(files) then iIn
         else if !isf.iovalue then deleteStaleDataFiles(isf.io, path, tail(files))
         else deleteStaleDataFiles( deleteFile(path ++ head(files), isf.io).io, path, tail(files));
}


