grammar silver:modification:autocopyattr;

build silver:modification:autocopyattr:java with silver:translation:java;

