grammar silver_construction;

imports silver:testing;

mainTestSuite silver_construction_tests;
