
imports lib:lsp;
imports lib:lsp:json;
