grammar silver:compiler:extension:monad;

imports silver:compiler:definition:core;
imports silver:compiler:definition:type:syntax;

imports silver:compiler:definition:env;
imports silver:compiler:definition:type;

imports silver:compiler:extension:convenience;
imports silver:compiler:modification:lambda_fn;
imports silver:compiler:modification:let_fix;

