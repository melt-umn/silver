grammar silver:modification:lambda_fn;

imports silver:definition:core;
imports silver:definition:env;
imports silver:definition:type;
imports silver:definition:type:syntax;
--imports silver:analysis:typechecking:core;

exports silver:modification:lambda_fn:java with silver:translation:java:core;
exports silver:modification:lambda_fn:java with silver:translation:java:type;

