grammar silver:host;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Host\nmenu_title: Host\nmenu_weight: 100\n---"
@}

