grammar tutorials:expr:host ;


import tutorials:expr:terminals ;
import tutorials:expr:abstractsyntax ;
import tutorials:expr:concretesyntax ;
import tutorials:expr:driver ;

