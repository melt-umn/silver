@@{-Docs in A.sv-}