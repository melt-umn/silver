grammar silver:core;

nonterminal Unit;

abstract production unit
top::Unit ::=
{}