grammar silver:compiler:modification:ffi;

exports silver:compiler:modification:ffi:java with silver:compiler:translation:java:core;

exports silver:compiler:modification:ffi:java with silver:compiler:translation:java:type;

