
imports lib:lsp;
imports core with deleteFile as COREdeleteFile;
