
-- annotation otxinfo :: OtxInfo;

-- nonterminal OtxInfo;
-- nonterminal OtxRule;
-- nonterminal OtxOriginLink;
