grammar silver:extension:autoattr;

terminal Propagate_kwd 'propagate' lexer classes {KEYWORD,RESERVED};
terminal Excluding_kwd 'excluding' lexer classes {KEYWORD};

terminal Functor_kwd   'functor' lexer classes {KEYWORD,RESERVED};
terminal Monoid_kwd    'monoid'  lexer classes {KEYWORD,RESERVED};
