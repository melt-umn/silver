grammar silver:core;

imports silver:core;
