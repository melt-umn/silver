grammar lib:lsp:document;

type DocumentUri = String;
synthesized attribute uri :: DocumentUri;
