grammar lib:monto:helpers;
