grammar test:nonterm_b_2;

nonterminal B;