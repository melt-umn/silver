
imports lib:lsp;
imports core with Location as CoreLocation;
