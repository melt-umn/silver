grammar silver:compiler:extension:abella_compilation:parsing_thms;

imports silver:compiler:extension:abella_compilation:abella;

--unparse attribute
imports silver:compiler:definition:core;

