import lib:json;

synthesized attribute json :: Json;
