grammar silver:extension:autoattr;

imports silver:definition:core;
imports silver:definition:env;
imports silver:definition:type;
imports silver:definition:type:syntax;
imports silver:modification:collection;
imports silver:modification:let_fix;
imports silver:extension:patternmatching;
imports silver:metatranslation;

exports silver:extension:autoattr:convenience;
