grammar silver:extension:constructparser;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Construct Parser\nmenu_title: Construct Parser\nmenu_weight: 100\n---"
@}

