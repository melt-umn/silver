grammar silver:compiler:modification:ffi;

{@config
  header:"---\nlayout: sv_wiki\ntitle: FFI\nmenu_title: FFI\nmenu_weight: 100\n---"
@}

