grammar silver:modification:collection;

exports silver:modification:collection:java with silver:translation:java;

