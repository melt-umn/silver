grammar silver:modification:collection:env_parser;

