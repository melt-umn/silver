grammar silver:compiler:modification:collection;

imports silver:compiler:definition:env;
imports silver:compiler:definition:core;
imports silver:compiler:definition:type;

exports silver:compiler:modification:collection:java with silver:compiler:translation:java:core;

