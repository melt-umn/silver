grammar silver_features:rewrite;

exports silver_features:rewrite:expreval;
