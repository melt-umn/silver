grammar silver:translation:java:command;

