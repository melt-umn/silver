grammar silver:compiler:extension:tuple;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Tuple\nmenu_title: Tuple\nmenu_weight: 100\n---"
@}