grammar lib:system ;

