imports doctest:split;
imports doctest:nonsplit;

@@{-@config excludeGrammar false-}