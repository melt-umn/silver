grammar lib;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Libraries\nmenu_title: Libraries\nmenu_weight: 100\n---"
@}

