grammar lib:lsp:hover;

imports lib:lsp;
imports lib:lsp:json;
imports lib:lsp:document;
