grammar silver:compiler:modification:collection;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Collections\nmenu_title: Collection\nmenu_weight: 100\n---"
@}

