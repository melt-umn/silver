
terminal Propagate_kwd 'propagate' lexer classes {KEYWORD,RESERVED};


