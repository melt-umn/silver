grammar silver:definition:core:env_parser;