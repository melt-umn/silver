grammar core;

synthesized attribute patProdName :: String;
synthesized attribute patChildList :: [AnyType];