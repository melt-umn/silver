grammar silver:xml:foreigntypes;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Foreign Types\nmenu_title: Foreign Types\nmenu_weight: 100\n---"
@}

