grammar silver:json;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Json\nmenu_title: Json\nmenu_weight: 100\n---"
@}

