grammar silver:compiler:modification:concisefunctions:java;

imports silver:compiler:definition:core;
imports silver:compiler:definition:env;
imports silver:compiler:definition:type;
imports silver:compiler:translation:java;
imports silver:compiler:analysis:typechecking:core;
imports silver:compiler:modification:concisefunctions;

