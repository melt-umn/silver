
annotation location :: Location;

