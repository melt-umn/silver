grammar silver_features:cond:e;

global cVal :: Integer = 9;

