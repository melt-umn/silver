grammar silver:modification:ffi;

build silver:modification:ffi:java with silver:translation:java;

