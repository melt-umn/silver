grammar silver:compiler:definition:core;

abstract production defaultAttributionDcl
top::AGDcl ::= at::Decorated QName attl::BracketedOptTypeExprs nt::QName nttl::BracketedOptTypeExprs
{
  top.unparse = "attribute " ++ at.unparse ++ attl.unparse ++ " occurs on " ++ nt.unparse ++ nttl.unparse ++ ";";

  -- TODO: this location is highly unreliable.

  -- We must unconditionally emit the occurs def in order to signal to the
  -- environment mechanism that we're in a different namespace than
  -- the types/attributes.
  top.occursDefs := [
    (if !at.lookupAttribute.dcl.isAnnotation then occursDcl else annoInstanceDcl)(
      nt.lookupType.fullName, at.lookupAttribute.fullName,
      protontty, protoatty,
      sourceGrammar=top.grammarName, sourceLocation=at.location)];

  -- binding errors in looking up these names.
  top.errors <- nt.lookupType.errors ++
    -- The nonterminal type list is strictly type VARIABLES only
    nttl.errorsTyVars;
  
  top.errors <-
    if attl.missingCount > 0
    then [err(attl.location, "Attribute type arguments cannot contain _")]
    else [];
  
  nttl.initialEnv = top.env;
  attl.env = nttl.envBindingTyVars;
  nttl.env = nttl.envBindingTyVars;
  
  local ntTypeScheme::PolyType = nt.lookupType.typeScheme;
  local atTypeScheme::PolyType = at.lookupAttribute.typeScheme;
  
  -- Make sure we get the number and kind of type variables correct for the NT
  top.errors <-
    case nt.lookupType.dcls of
    | ntDcl(_, ks, _, _) :: _ when length(ks) != length(nttl.types) ->
      [err(nt.location,
        nt.name ++ " expects " ++ toString(length(ks)) ++
        " type variables, but " ++ toString(length(nttl.types)) ++ " were provided.")]
    | ntDcl(_, ks, _, _) :: _ when ks != map((.kindrep), nttl.types) ->
      [err(nt.location,
        nt.name ++ " had kind " ++ foldr(arrowKind, starKind(), ks).typepp ++
        "but type variable(s) have kind(s) " ++ implode(", ", map(compose(prettyKind, (.kindrep)), nttl.types)) ++ ".")]
    | _ -> []
    end;

  -- Make sure we get the number and kind of type variables correct for the ATTR
  top.errors <-
    if length(atTypeScheme.boundVars) != length(attl.types)
    then [err(at.location,
      at.name ++ " expects " ++ toString(length(atTypeScheme.boundVars)) ++
      " type variables, but " ++ toString(length(attl.types)) ++ " were provided.")]
    else if map((.kindrep), atTypeScheme.boundVars) != map((.kindrep), attl.types)
    then [err(at.location,
      at.name ++ " has kind " ++ prettyKind(foldr(arrowKind, starKind(), map((.kindrep), atTypeScheme.boundVars))) ++
        "but type variable(s) have kind(s) " ++ implode(", ", map(compose(prettyKind, (.kindrep)), attl.types)) ++ ".")]
    else [];

  -- We have 4 types.
  -- 1: A type, from env, for the nonterminal (unapplied)
  -- 2: A type, from syntax, for the nonterminal (applied to type vars)
  -- 3: A type, from env, for the attribute (with bound type vars)
  -- 4: A type, from syntax, for the attribute (sharing the same type vars as #2)
  
  -- Our goal is to be able to take a (unknown) nonterminal type
  -- and yield the appropriate attribute type it corresponds to.
  
  -- To that end, we want two things:
  -- 1: A type that we can unify with some nonterminal type.
  -- 2: A type that, under that unification, will be the resulting attribute type.

  -- So we generate a list of fresh type variables corresponding to the types of #2,
  -- and generate two substitutions:
  -- 1: Rewrite the tyvars of type #3 to the types of type #4.
  -- 2: Rewrite our local tyvars to fresh variables.
  
  -- Thus, we apply #1 to our fresh type vars, perform both substitutions on #3, and get our goal.
  
  -- Fresh type variables that will go in the environment
  local tyVars :: [TyVar] = freshTyVars(nttl.freeVariables);
  
  -- Apply the nonterminal type to the type variables.
  -- NOT .monoType so we do something sensible if someone does "occurs on TypeAlias<a>" or something.
  production protontty :: Type = appTypes(ntTypeScheme.typerep, map(varType, tyVars));
  
  -- This renames the vars from the environment
  -- at's env types -> type params containing local skolem vars  (vars -> types)
  local rewrite_from :: Substitution = zipVarsAndTypesIntoSubstitution(atTypeScheme.boundVars, attl.types);
  
  -- local skolem vars -> fresh type vars (vars -> vars)
  local rewrite_to :: Substitution = zipVarsIntoSubstitution(nttl.freeVariables, tyVars);
  
  -- These have to be two separate renamings, because the second renaming replaces names getting substituted in by the first renaming.
  production protoatty :: Type = performRenaming(performRenaming(atTypeScheme.typerep, rewrite_from), rewrite_to);
  
  -- Now, finally, make sure we're not "redefining" the occurs.
  production occursCheck :: [DclInfo] = getOccursDcl(at.lookupAttribute.fullName, nt.lookupType.fullName, top.env);
  
  top.errors <-
    if length(occursCheck) > 1
    then [err(at.location, "Attribute '" ++ at.name ++ "' already occurs on '" ++ nt.name ++ "'.")]
    else [];

  top.errors <-
    if nt.lookupType.found && (!nt.lookupType.dcl.isType || !ntTypeScheme.typerep.isDecorable)
    then [err(nt.location, nt.name ++ " is not a nonterminal. Attributes can only occur on nonterminals.")]
    else [];
                
  top.errors <-
    if !nt.lookupType.found || !at.lookupAttribute.found || !at.lookupAttribute.dcl.isAnnotation ||
       isExportedBy(top.grammarName, [nt.lookupType.dcl.sourceGrammar], top.compiledGrammars) then []
    else [err(top.location, "Annotations for a nonterminal must be in a module exported by the nonterminal's declaring grammar.")];
}

abstract production errorAttributionDcl
top::AGDcl ::= msg::[Message] at::Decorated QName attl::BracketedOptTypeExprs nt::QName nttl::BracketedOptTypeExprs
{
  top.unparse = "attribute " ++ at.unparse ++ attl.unparse ++ " occurs on " ++ nt.unparse ++ nttl.unparse ++ ";";
  top.occursDefs := [];
  top.errors <- msg;
  
  nttl.initialEnv = top.env;
  attl.env = nttl.envBindingTyVars;
  nttl.env = nttl.envBindingTyVars;
  
  -- Decorate everything else to still check for errors
  top.errors <-
    -- binding errors in looking up these names.
    nt.lookupType.errors ++
    -- The nonterminal type list is strictly type VARIABLES only
    nttl.errorsTyVars;
  
  -- Make sure we get the number and kinds of tyvars correct for the NT
  top.errors <-
    case nt.lookupType.dcls of
    | ntDcl(_, ks, _, _) :: _ when length(ks) != length(nttl.types) ->
      [err(nt.location,
        nt.name ++ " expects " ++ toString(length(ks)) ++
        " type variables, but " ++ toString(length(nttl.types)) ++ " were provided.")]
    | ntDcl(_, ks, _, _) :: _ when ks != map((.kindrep), nttl.types) ->
      [err(nt.location,
        nt.name ++ " had kind " ++ foldr(arrowKind, starKind(), ks).typepp ++
        "but type variable(s) have kind(s) " ++ implode(", ", map(compose(prettyKind, (.kindrep)), nttl.types)) ++ ".")]
    | _ -> []
    end;
}

concrete production attributionDcl
top::AGDcl ::= 'attribute' at::QName attl::BracketedOptTypeExprs 'occurs' 'on' nt::QName nttl::BracketedOptTypeExprs ';'
{
  top.unparse = "attribute " ++ at.unparse ++ attl.unparse ++ " occurs on " ++ nt.unparse ++ nttl.unparse ++ ";";
  
  -- Workaround for circular dependency due to dispatching on env:
  -- Nothing used to build the env namespaces on which we dispatch can depend on
  -- the forward here.
  -- Attribution (occurs) defs, which obviously must depend on this forward, are
  -- specified by a separate occursDefs attribute.
  -- Attribution dispatch productions should only define occursDefs (i.e. no new
  -- nonterminals, productions, attributes, etc.)
  top.defs := [];
  top.moduleNames := [];
  
  forwards to
    (if !at.lookupAttribute.found
     then errorAttributionDcl(at.lookupAttribute.errors, _, _, _, _, location=_)
     else at.lookupAttribute.dcl.attributionDispatcher)(at, attl, nt, nttl, top.location);
}

concrete production annotateDcl
top::AGDcl ::= 'annotation' at::QName attl::BracketedOptTypeExprs 'occurs' 'on' nt::QName nttl::BracketedOptTypeExprs ';'
{
  forwards to attributionDcl('attribute', at, attl, $4, $5, nt, nttl, $8, location=top.location);
}

