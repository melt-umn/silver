grammar core;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Core library\nmenu_title: core library\nmenu_weight: 20\n---"

  split-files: "true"
@}

