grammar tutorial:expr:terminals ;

terminal Fst_t     'fst' dominates { Id_t } ;
terminal Snd_t     'snd' dominates { Id_t } ;

