grammar silver:modification:copper;

imports silver:definition:core;
imports silver:definition:env;
imports silver:definition:concrete_syntax;
imports silver:definition:concrete_syntax:ast;
imports silver:definition:type;
imports silver:definition:type:syntax;

imports silver:analysis:typechecking:core;
imports silver:analysis:typechecking;

imports silver:translation:java:core;
imports silver:translation:java:type;

imports silver:util;

