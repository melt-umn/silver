@@{-Doc-}