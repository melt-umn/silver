
terminal Propagate_kwd 'propagate' lexer classes {KEYWORD,RESERVED};
terminal Functor_kwd   'functor' lexer classes {KEYWORD,RESERVED};
