grammar core;

imports core:monad;
imports core:reflect;
