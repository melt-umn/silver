grammar silver_features ;

imports silver:testing ;
imports lib:extcore ;

mainTestSuite silver_tests ;

