grammar silver:compiler:modification:lambda_fn;

{@config
  header:"---\nlayout: sv_wiki\ntitle: Lambda Functions\nmenu_title: Lambda Functions\nmenu_weight: 100\n---"
@}

