
terminal Propagate_kwd 'propagate' lexer classes {KEYWORD,RESERVED};
terminal PropagateOld_kwd 'propagate_functor' lexer classes {KEYWORD,RESERVED};
terminal Functor_kwd   'functor' lexer classes {KEYWORD,RESERVED};
