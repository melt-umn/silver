function nutshack
Integer ::= {return 0;}