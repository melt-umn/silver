grammar tutorials:expr:terminals ;


terminal Input_t  'input' dominates { Id_t } ;

terminal Comma_t    ','  ;
