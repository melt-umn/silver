grammar silver:analysis:typechecking:type:io;
export silver:analysis:typechecking:type:io;
