grammar silver:core;

@@{-
   - @config split
   - @config grammarWeight -1
   - @config grammarTitle "[silver:core] (stdlib)"
   -}