grammar silver:extension:templating;

{@config
  header:"---\nlayout: sv_wiki\ntitle: String Templating\nmenu_title: String Templating\nmenu_weight: 100\n---"
@}

